//Add
module add(a1,a2,yout);
input [27:0]a1;
input [31:0]a2;
output [31:0]yout;
assign yout=a1+a2;
endmodule
