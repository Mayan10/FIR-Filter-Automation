//Adder21
module adder21(a,b,c  );
input [31:0]a;
input [39:0]b;
output  [39:0]c;
assign c=a+b;
endmodule
