
//Adder22
module adder22(a,b,c  );
input [39:0]a;
input [47:0]b;
output [47:0]c;
assign c=a+b;
endmodule
