//Adder
module adder(a,b,c);
input [27:0]a;
input [27:0]b;
output  [27:0]c;
assign c=a+b;
endmodule
